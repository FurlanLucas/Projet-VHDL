library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity windowing_TB is
end entity;

architecture windowing_TB_arch of windowing_TB is

	component windowing
		port(CLK    : in std_logic;
		     CE     : in std_logic;
			 reset  : in std_logic;
			 entree : in std_logic_vector(11 downto 0);
			 sortie: out std_logic_vector(11 downto 0);
			 test : out std_logic);
	end component;
	
	signal CLK_TB    : std_logic;
	signal CE_TB     : std_logic;
	signal reset_TB  : std_logic;
 	signal entree_TB : std_logic_vector(11 downto 0);
	signal sortie_TB : std_logic_vector(11 downto 0);
	signal test_TB :  std_logic;
	
begin

	DUT : windowing port map(CLK => CLK_TB,
	                            CE => CE_TB,
								reset => reset_TB,
								entree => entree_TB,
								sortie => sortie_TB,
								test => test_TB);
				
	CLK : process
	begin
		CLK_TB <= '1';
		wait for 5 ns;
		CLK_TB <= '0';
		wait for 5 ns;
	end process;
	
    CE : process
	begin
		CE_TB <= '0';
		wait for 390 ns;
		CE_TB <= '1';
		wait for 10 ns;
	end process;

	RST : process
	begin
		reset_TB <= '1';
		wait for 10 ns;
		reset_TB <= '0';
		wait for 100 ms;
	end process;
	
	SMT : process
	begin
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011001000";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000111";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000110";
        wait for 400 ns;
        entree_TB <= "000011000101";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000100";
        wait for 400 ns;
        entree_TB <= "000011000011";
        wait for 400 ns;
        entree_TB <= "000011000010";
        wait for 400 ns;
        entree_TB <= "000011000001";
        wait for 400 ns;
        entree_TB <= "000010111111";
        wait for 400 ns;
        entree_TB <= "000010111110";
        wait for 400 ns;
        entree_TB <= "000010111101";
        wait for 400 ns;
        entree_TB <= "000010111011";
        wait for 400 ns;
        entree_TB <= "000010111010";
        wait for 400 ns;
        entree_TB <= "000010111000";
        wait for 400 ns;
        entree_TB <= "000010110111";
        wait for 400 ns;
        entree_TB <= "000010110101";
        wait for 400 ns;
        entree_TB <= "000010110011";
        wait for 400 ns;
        entree_TB <= "000010110001";
        wait for 400 ns;
        entree_TB <= "000010101111";
        wait for 400 ns;
        entree_TB <= "000010101101";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000000000";
        wait for 400 ns;
        entree_TB <= "000000000100";
        wait for 400 ns;
        entree_TB <= "000000001000";
        wait for 400 ns;
        entree_TB <= "000000001101";
        wait for 400 ns;
        entree_TB <= "000000010001";
        wait for 400 ns;
        entree_TB <= "000000010101";
        wait for 400 ns;
        entree_TB <= "000000011001";
        wait for 400 ns;
        entree_TB <= "000000011101";
        wait for 400 ns;
        entree_TB <= "000000100001";
        wait for 400 ns;
        entree_TB <= "000000100101";
        wait for 400 ns;
        entree_TB <= "000000101010";
        wait for 400 ns;
        entree_TB <= "000000101110";
        wait for 400 ns;
        entree_TB <= "000000110010";
        wait for 400 ns;
        entree_TB <= "000000110110";
        wait for 400 ns;
        entree_TB <= "000000111010";
        wait for 400 ns;
        entree_TB <= "000000111110";
        wait for 400 ns;
        entree_TB <= "000001000010";
        wait for 400 ns;
        entree_TB <= "000001000110";
        wait for 400 ns;
        entree_TB <= "000001001010";
        wait for 400 ns;
        entree_TB <= "000001001110";
        wait for 400 ns;
        entree_TB <= "000001010001";
        wait for 400 ns;
        entree_TB <= "000001010101";
        wait for 400 ns;
        entree_TB <= "000001011001";
        wait for 400 ns;
        entree_TB <= "000001011101";
        wait for 400 ns;
        entree_TB <= "000001100000";
        wait for 400 ns;
        entree_TB <= "000001100100";
        wait for 400 ns;
        entree_TB <= "000001101000";
        wait for 400 ns;
        entree_TB <= "000001101011";
        wait for 400 ns;
        entree_TB <= "000001101111";
        wait for 400 ns;
        entree_TB <= "000001110010";
        wait for 400 ns;
        entree_TB <= "000001110110";
        wait for 400 ns;
        entree_TB <= "000001111001";
        wait for 400 ns;
        entree_TB <= "000001111100";
        wait for 400 ns;
        entree_TB <= "000001111111";
        wait for 400 ns;
        entree_TB <= "000010000011";
        wait for 400 ns;
        entree_TB <= "000010000110";
        wait for 400 ns;
        entree_TB <= "000010001001";
        wait for 400 ns;
        entree_TB <= "000010001100";
        wait for 400 ns;
        entree_TB <= "000010001111";
        wait for 400 ns;
        entree_TB <= "000010010010";
        wait for 400 ns;
        entree_TB <= "000010010101";
        wait for 400 ns;
        entree_TB <= "000010010111";
        wait for 400 ns;
        entree_TB <= "000010011010";
        wait for 400 ns;
        entree_TB <= "000010011101";
        wait for 400 ns;
        entree_TB <= "000010011111";
        wait for 400 ns;
        entree_TB <= "000010100010";
        wait for 400 ns;
        entree_TB <= "000010100100";
        wait for 400 ns;
        entree_TB <= "000010100111";
        wait for 400 ns;
        entree_TB <= "000010101001";
        wait for 400 ns;
        entree_TB <= "000010101011";
        wait for 400 ns;

		
	end process;
	
end architecture;